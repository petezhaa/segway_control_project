module Segway_tb ();

  import task_pkg::*;

  //// Interconnects to DUT/support defined as type wire /////
  wire SS_n, SCLK, MOSI, MISO, INT;  // to inertial sensor
  wire A2D_SS_n, A2D_SCLK, A2D_MOSI, A2D_MISO;  // to A2D converter
  wire RX_TX;
  wire PWM1_rght, PWM2_rght, PWM1_lft, PWM2_lft;
  wire piezo, piezo_n;
  wire cmd_sent;
  wire rst_n;  // synchronized global reset

  ////// Stimulus is declared as type reg ///////
  reg clk, RST_n;
  reg [7:0] cmd;  // command host is sending to DUT
  reg send_cmd;  // asserted to initiate sending of command
  reg signed [15:0] rider_lean;
  reg [11:0] ld_cell_lft, ld_cell_rght, steerPot, batt;  // A2D values
  reg OVR_I_lft, OVR_I_rght;

  ///// Internal registers for testing purposes??? /////////

  ////////////////////////////////////////////////////////////////
  // Instantiate Physical Model of Segway with Inertial sensor //
  //////////////////////////////////////////////////////////////	
  SegwayModel iPHYS (
      .clk(clk),
      .RST_n(RST_n),
      .SS_n(SS_n),
      .SCLK(SCLK),
      .MISO(MISO),
      .MOSI(MOSI),
      .INT(INT),
      .PWM1_lft(PWM1_lft),
      .PWM2_lft(PWM2_lft),
      .PWM1_rght(PWM1_rght),
      .PWM2_rght(PWM2_rght),
      .rider_lean(rider_lean)
  );

  /////////////////////////////////////////////////////////
  // Instantiate Model of A2D for load cell and battery //
  ///////////////////////////////////////////////////////
  ADC128S_FC iA2D (
      .clk(clk),
      .rst_n(RST_n),
      .SS_n(A2D_SS_n),
      .SCLK(A2D_SCLK),
      .MISO(A2D_MISO),
      .MOSI(A2D_MOSI),
      .ld_cell_lft(ld_cell_lft),
      .ld_cell_rght(ld_cell_rght),
      .steerPot(steerPot),
      .batt(batt)
  );

  ////// Instantiate DUT ////////
  Segway iDUT (
      .clk(clk),
      .RST_n(RST_n),
      .INERT_SS_n(SS_n),
      .INERT_MOSI(MOSI),
      .INERT_SCLK(SCLK),
      .INERT_MISO(MISO),
      .INERT_INT(INT),
      .A2D_SS_n(A2D_SS_n),
      .A2D_MOSI(A2D_MOSI),
      .A2D_SCLK(A2D_SCLK),
      .A2D_MISO(A2D_MISO),
      .PWM1_lft(PWM1_lft),
      .PWM2_lft(PWM2_lft),
      .PWM1_rght(PWM1_rght),
      .PWM2_rght(PWM2_rght),
      .OVR_I_lft(OVR_I_lft),
      .OVR_I_rght(OVR_I_rght),
      .piezo_n(piezo_n),
      .piezo(piezo),
      .RX(RX_TX)
  );

  //// Instantiate UART_tx (mimics command from BLE module) //////
  UART_tx iTX (
      .clk(clk),
      .rst_n(rst_n),
      .TX(RX_TX),
      .trmt(send_cmd),
      .tx_data(cmd),
      .tx_done(cmd_sent)
  );

  /////////////////////////////////////
  // Instantiate reset synchronizer //
  ///////////////////////////////////
  rst_synch iRST (
      .clk  (clk),
      .RST_n(RST_n),
      .rst_n(rst_n)
  );

  initial begin

    /// Your magic goes here /// // use connect by name here 
    init_DUT(.clk(clk), .RST_n(RST_n), .send_cmd(send_cmd), .cmd(cmd), .rider_lean(rider_lean),
             .ld_cell_lft(ld_cell_lft), .ld_cell_rght(ld_cell_rght), .steerPot(steerPot),
             .batt(batt), .OVR_I_lft(OVR_I_lft), .OVR_I_rght(OVR_I_rght));

    // Send 'G' command
    SendCmd(.clk(clk), .trmt(send_cmd), .tx_data(cmd), .cmd(G));

    ld_cell_lft  = 12'h300;  // simulate rider getting on
    ld_cell_rght = 12'h300;  // simulate rider getting on
    repeat (350000) @(posedge clk);  // wait for some time

    rider_lean = 16'sh0FFF;  // simulate rider leaning forward

    repeat (1000000) @(posedge clk);  // wait for some time

    // ----------------------------------------------------------
    // 5) Abruptly remove lean (back to zero) and watch ring-down
    // ----------------------------------------------------------
    rider_lean = 16'sh0000;
    repeat (800000) @(posedge clk);  // wait for some time


    // ================== Added Comprehensive System Tests ==================

    // Steering right then left (differential wheel response)
    steerPot = 12'hE00;
    repeat (600000) @(posedge clk);
    steerPot = 12'h200;
    repeat (600000) @(posedge clk);
    steerPot = 12'h800; // center
    repeat (300000) @(posedge clk);

    // Rider lean forward then backward (speed reversal / braking)
    rider_lean = 16'sh0600;
    repeat (800000) @(posedge clk);
    rider_lean = -16'sh0400;
    repeat (800000) @(posedge clk);
    rider_lean = 16'sh0000;
    repeat (400000) @(posedge clk);

    // Simulate step-off (load cells go low) -> expect internal disable
    ld_cell_lft  = 12'h020;
    ld_cell_rght = 12'h010;
    repeat (600000) @(posedge clk);

    // Re-mount rider and send STOP then GO sequence
    ld_cell_lft  = 12'h300;
    ld_cell_rght = 12'h300;
    repeat (200000) @(posedge clk);
    SendCmd(.clk(clk), .trmt(send_cmd), .tx_data(cmd), .cmd(S));
    repeat (400000) @(posedge clk);
    SendCmd(.clk(clk), .trmt(send_cmd), .tx_data(cmd), .cmd(G));
    repeat (600000) @(posedge clk);

    // Transient overcurrent pulse (left)
    OVR_I_lft = 1;
    repeat (2000) @(posedge clk);
    OVR_I_lft = 0;
    repeat (300000) @(posedge clk);

    // Persistent overcurrent (right)
    OVR_I_rght = 1;
    repeat (1_200_000) @(posedge clk);
    OVR_I_rght = 0;
    repeat (300000) @(posedge clk);

    // Dual overcurrent short event
    OVR_I_lft  = 1;
    OVR_I_rght = 1;
    repeat (300000) @(posedge clk);
    OVR_I_lft  = 0;
    OVR_I_rght = 0;
    repeat (300000) @(posedge clk);

    // Battery voltage ramp down (warning / shutdown behavior)
    batt = 12'hC00;
    repeat (200000) @(posedge clk);
    batt = 12'hA00;
    repeat (200000) @(posedge clk);
    batt = 12'h800;
    repeat (200000) @(posedge clk);
    batt = 12'h650;
    repeat (300000) @(posedge clk);
    batt = 12'h500; // near critical
    repeat (400000) @(posedge clk);
    batt = 12'h3A0; // critical low
    repeat (400000) @(posedge clk);

    // Simulate fall (excessive tilt)
    rider_lean = 16'sh1FFF;
    repeat (600000) @(posedge clk);
    rider_lean = 16'sh0000;
    repeat (400000) @(posedge clk);

    // Final STOP
    SendCmd(.clk(clk), .trmt(send_cmd), .tx_data(cmd), .cmd(S));
    repeat (400000) @(posedge clk);

    // ======================================================================

    #100;
    $stop();
  end

  always #10 clk = ~clk;

endmodule